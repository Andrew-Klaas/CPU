module cache_datapath
(
   input    logic          clk,
   
   // Cache Datapath <--> CPU
   input    logic[1:0]     mem_byte_enable,
   input    logic[15:0]    mem_address,
   input    logic[15:0]    mem_wdata,
   input    logic          mem_write,
   output   logic[15:0]    mem_rdata,
   
   // Cache Datapath <--> Cache Control
   input    logic          L_in,
   input    logic          WE0,
   input    logic          WE1,
   input    logic          WEL,
   input    logic          D0_in,
   input    logic          D1_in,
   input    logic          feedback_sel,
   input    logic          output_mode,
   input    logic          output_set,
   output   logic          hit,
   output   logic          hit_set,
   output   logic          V0_out,
   output   logic          V1_out,
   output   logic          D0_out,
   output   logic          D1_out,
   output   logic          L_out,
   
   // Cache Datapath <--> Physical Memory
   input    logic[127:0]   pmem_rdata,
   output   logic[127:0]   pmem_wdata,
   output   logic[15:0]    pmem_address,
   
   // peeking circuitry added to support prefetching
   input    logic[15:0]    peek_address,
   output   logic          peek_hit
   
);
   
   /* Instantiate the actual cache lines
    * Since this is a 2-way set associative cache, there will be two ways.
    * Each way has 8 cache lines, selected using ix == mem_address[5:3].
    * Each of these lines has a valid bit (V), 10-bit tag (mem_address[15:6])
    * and a 128-bit cache line. Data is written to all 3 elements at once
    * whenever WE == 1 during a rising clock edge */
   
   logic[127:0]      data0_out;
   logic[8:0]        tag0_out;
   
   logic[127:0]      data1_out;
   logic[8:0]        tag1_out;
   
   logic[127:0]      merge_out;
   
   logic             peek_hit0;
   logic             peek_hit1;
   
   cache_way   WAY0_INST
   (
      .clk,
      .WE(WE0),
      .ix(mem_address[6:4]),
      
      .D_in(D0_in),
      .tag_in(mem_address[15:7]),
      .data_in(merge_out),
      
      .V_out(V0_out),
      .D_out(D0_out),
      .tag_out(tag0_out),
      .data_out(data0_out),
      
      .peek_address,
      .peek_hit(peek_hit0)
   );
   
   cache_way   WAY1_INST
   (
      .clk,
      .WE(WE1),
      .ix(mem_address[6:4]),
      
      .D_in(D1_in),
      .tag_in(mem_address[15:7]),
      .data_in(merge_out),
      
      .D_out(D1_out),
      .V_out(V1_out),
      .tag_out(tag1_out),
      .data_out(data1_out),
      
      .peek_address,
      .peek_hit(peek_hit1)
   );
   
   assign   peek_hit = peek_hit0 || peek_hit1;
   
   L_array L_ARRAY_INST
   (
      .clk,
      .WE(WEL),
      .ix(mem_address[6:4]),
      .L_in,
      .L_out
   );
   
   /* The following code is two layers of multiplexers.
    * The first multiplexer is a 2-input, 128-bit MUX which
    * selects the data output from either way0 or way1 based
    * on the 'output_set' input pin.  The second MUX is an
    * 8-input,16-bit mux which selects one of the 16-bit words
    * out of the cache line and presents it to the CPU */
   always_comb
   begin
      
      // first multiplexer.  This selects the cache line from way0 or way1
      pmem_wdata = output_set ? data1_out : data0_out;
      
      // second multiplexer.  This selects a 16-bit word for the CPU
      case (mem_address[3:1])
         // even addresses only
         3'b000:     mem_rdata = pmem_wdata[15:0];
         3'b001:     mem_rdata = pmem_wdata[31:16];
         3'b010:     mem_rdata = pmem_wdata[47:32];
         3'b011:     mem_rdata = pmem_wdata[63:48];
         3'b100:     mem_rdata = pmem_wdata[79:64];
         3'b101:     mem_rdata = pmem_wdata[95:80];
         3'b110:     mem_rdata = pmem_wdata[111:96];
         3'b111:     mem_rdata = pmem_wdata[127:112];
         endcase
   end
   
   /* Caclulate the hit and hit_set bits */
   assign   hit_set  =  V1_out && (mem_address[15:7] == tag1_out);
   assign   hit      = (V0_out && (mem_address[15:7] == tag0_out)) || hit_set;
   
   /* Calculate the physical address.
    * If an eviction is is progress, then the tag from the evicted
    * cache line is gated to the physical address output.
    * If a fetch is in progress, then the address generated by the
    * CPU is gated to the physical address output */
   assign   pmem_address[15:7] = output_mode ? (output_set ? tag1_out : tag0_out) : mem_address[15:7]; // Tag
   assign   pmem_address[6:0]  = mem_address[6:0];  // Index.  The low 4 bits don't matter
   
   /* Circuitry for writing data from mem_wdata into a cache line */
   write_merge WRITE_MERGE_INST
   (
      .mem_write,
      .mem_byte_enable,
      .word_sel(mem_address[3:1]),
      
      .mem_wdata,
      .cache_line_in(feedback_sel ? pmem_wdata : pmem_rdata),
      .cache_line_out(merge_out)
   );
   
endmodule : cache_datapath
